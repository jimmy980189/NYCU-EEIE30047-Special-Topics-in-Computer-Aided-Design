module           
c17 (N1, 
    N2, 


    N3, N6, N7, N22, N23);
     
   wire n8, 
       n9, 
       n10, n11, n12;
	input
    N1, N2, N3, N6, N7;
 
	output /*adasd*//*dasd*/ N22, N/*;*/23; /*N24
// asdsadsad sadsadsadsadsad
    NOR2X1      
    U8 (./*.A0(fucku*/A1(n8),   .A2(n9),  /*A2(n8)
    */.ZN(N23));
	  NOR2X1 U9 (.A1(N2), /*sadsadas*/.A2(N7), .ZN(n9));//dhjikb/*
	INVX1 U10 (.I(n10), /*AAAAdsadsadsad*/ .ZN(n8));   //dgbou/*missme?*/
    // dasdsadsadsad 
            NANDX1 U11 (.A1(n11), .A2(n12),
             .ZN(N22)); //dsadsadsdsadsad
	NANDX1                   U12 (.A1(N2),   /*aaasdsad*/ .A2(n10), .ZN(n12))/* dsfdsfdsfjhhjhkjhjhd NANDX1 U11 (.A1(n11), .A2(n12), /* */;
	    /*asdsadsadsadasdsadsa*/NANDX1 U13 (.A1(N6),
          .A2(N3), .ZN(n10));
	NANDX1              U14    (.A1(N1), .A2(N3), /*sadsadsadasdasd*/.ZN(n11));
endmodule










